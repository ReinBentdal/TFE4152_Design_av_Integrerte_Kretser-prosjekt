
`ifndef _PIXEL_SENSOR_CONFIG
`define _PIXEL_SENSOR_CONFIG
package PixelSensorConfig;

    parameter PIXEL_ARRAY_HEIGHT = 2;
    parameter PIXEL_ARRAY_WIDTH = 2;

    parameter OUTPUT_BUS_WIDTH = 64;
endpackage
`endif