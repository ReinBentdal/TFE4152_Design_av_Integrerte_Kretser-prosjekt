

module readout();

    parameter bus_width = 64;    

endmodule