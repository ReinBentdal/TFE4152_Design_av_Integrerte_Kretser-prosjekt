`include "../../pixel_sensor_config.sv"

module readout(
    
    output data_out,
    output data_out_clk
);



    parameter bus_width = 64;



endmodule